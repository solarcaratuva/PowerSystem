*---------- DMP2110UW Spice Model ----------
.SUBCKT DMP2110UW 10 20 30 
*     TERMINALS:  D  G  S
M1 1 2 3 3 PMOS L = 1E-006 W = 1E-006 
RD 10 1 0.04439 
RS 30 3 0.001 
RG 20 2 8.47 
CGS 2 3 3.947E-010 
EGD 12 30 2 1 1 
VFB 14 30 0 
FFB 2 1 VFB 1 
CGD 13 14 7.7E-010 
R1 13 30 1 
D1 13 12 DLIM 
DDG 14 15 DCGD 
R2 12 15 1 
D2 30 15 DLIM 
DSD 10 3 DSUB 
.MODEL PMOS PMOS LEVEL = 3 U0 = 400 VMAX = 1E+006 ETA = 0.001 
+ TOX = 6E-008 NSUB = 1E+016 KP = 28.79 KAPPA = 19.32 VTO = -0.919 
.MODEL DCGD D CJO = 4.315E-010 VJ = 0.6 M = 0.7569 
.MODEL DSUB D IS = 1.86E-008 N = 1.276 RS = 0.06967 BV = 27 CJO = 7.361E-011 VJ = 0.6 M = 0.6276 TT = 4.2E-009 
.MODEL DLIM D IS = 0.0001 
.ENDS
*Diodes DMP2110UW Spice Model v1.0M Last Revised 2018/2/2